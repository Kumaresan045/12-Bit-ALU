module and81 (input [7:0] op1,input op2, output [7:0] out);

    and andi[7:0] (out[7:0],op1[7:0],op2);

endmodule