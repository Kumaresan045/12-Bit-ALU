module and41 (input [3:0] op1,input op2, output [3:0] out);

    and andi[3:0] (out[3:0],op1[3:0],op2);

endmodule