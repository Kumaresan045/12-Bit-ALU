module fa(input a, input b,input cin,output s,output cout);

    ha ha1 (a,b,p,g);
    ha ha2 (p,cin,s,temp);
    or (cout,g,temp);

endmodule