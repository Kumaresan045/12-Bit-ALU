module and12_1 (input [11:0] op1,input op2, output [11:0] out);

    and andi[11:0] (out[11:0],op1[11:0],op2);

endmodule