module and71 (input [6:0] op1,input op2, output [6:0] out);

    and andi[6:0] (out[6:0],op1[6:0],op2);

endmodule